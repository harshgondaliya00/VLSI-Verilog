`timescale 1ns / 1ps

module mux_tb;
    reg [3:0] s;
    reg [15:0] d;
    wire y;
    
    mux uut (
        .y(y),
        .s(s),
        .d(d)
    );

    initial begin
       
        s = 4'b0000; d = 16'h0001; #10; 
        s = 4'b0001; d = 16'h0002; #10;
        s = 4'b0010; d = 16'h0004; #10;
        s = 4'b0011; d = 16'h0008; #10;
        s = 4'b0100; d = 16'h0010; #10;
        s = 4'b0101; d = 16'h0020; #10;
        s = 4'b0110; d = 16'h0040; #10;
        s = 4'b0111; d = 16'h0080; #10;
        s = 4'b1000; d = 16'h0100; #10;
        s = 4'b1001; d = 16'h0200; #10;
        s = 4'b1010; d = 16'h0400; #10;
        s = 4'b1011; d = 16'h0800; #10;
        s = 4'b1100; d = 16'h1000; #10;
        s = 4'b1101; d = 16'h2000; #10;
        s = 4'b1110; d = 16'h4000; #10;
        s = 4'b1111; d = 16'h8000; #10;


        $finish;
    end
endmodule
